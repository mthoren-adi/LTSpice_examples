
.subckt CUSTOMBLOCK 1 2 3 4 5 6 7
CG1 117 0 2.9E-7
CG3 118 0 5E-7
CIN1 3 2 4p
CIN2 2 4 4p
CIN3 3 5 4p
CIN4 5 4 4p
CPSRR1 114 119 1.2p
DIN1 5 112 DIN
DIN2 112 113 DIN
DIN3 113 22 DIN
DIN4 21 22 DIN
DIN5 22 21 DIN
DVL1 116 117 DVLIM1
DVL2 116 0 DVLIM2
DZ1 3 5 DZNR
DZ2 2 1 DZNR
EVLIM1 119 0 5 0 1
EVLIM2 120 0 VALUE={V(5)-4}
GG1 0 117 VALUE={4*TANH(V(23))}
GG3 0 118 117 0 6.2832
GGAIN 0 23 111 22 1.5625m
GINX1 0 111 21 0 1
GOUT 0 121 118 0 10m
GPSRR 0 122 5 2 5.62e-12
GPSRRO 111 0 122 0 1
GPWR 5 2 115 0 1E-6
IBIAS1 21 0 1.5n
IBIAS2 22 0 1.5n
IOS 21 22 2n
ISUPTC 0 115 1
IVOS 0 111 20u
MCUR 1a 6a 6 6 PCUR
*MCUR 1 6a 6 6 PCUR
MOUT1 119 121 6a 6a NOUT
MOUT2 120 121 6a 6a POUT
RA 23 0 800
RG1 117 0 160K
RG3 118 0 0.159155
RIN1 21 4 5k
RIN2 22 3 5k
RINX1 111 0 1
ROUT1 119 121 200
ROUT2 121 120 200
RPSRR1 122 0 1k
RPSRR2 122 114 1meg
RPWR 2 5 440k
RSUPTC 115 0 210 TC1=5m

* SHDN
* SHDN pin has ESD (DZ3)
* SHDN pin has Series 5K (RSHDN)
* Protection after 5K (DVL7)
* Inverter (M11 and M12)
* Output pass transistor (MCUTOFF)
* Protection for MCUTOFF drain (DZ4)
* MCUTOFF bridges main circuit 1a to output 1
* 5 V supply V5V acts to do what proper circuitry would
* do, namely keep a small supply alive to run the inverter logic.
DZ3 2 7 DZNR
DVL7 2 140 DZNR
DZ4 2 1a DZNR
M11 142 140 141 141 PMOSGEN
M12 142 140 2 2 NMOSGEN
MCUTOFF 1a 142 1 1 NCUR
RSHDN 7 140 5K
RSIM 1a 1 1000Meg
V5V 141 2 DC 5


.MODEL NCUR NMOS(KF=0 KP=5E-4)

.MODEL NOUT NMOS(KF=0 KP=5 VTO=-10M)
.MODEL POUT PMOS(KF=0 KP=5 VTO=10M)
.MODEL PCUR PMOS(KF=0 KP=5E-4)
.MODEL NMOSGEN NMOS
.MODEL PMOSGEN PMOS
.MODEL DIN D(KF=0 RS=0)
.MODEL DVLIM1 D(BV=1.2 IS=1E-10 KF=0 RS=0)
.MODEL DVLIM2 D(BV=5 IS=1E-10 KF=0 RS=0)
.MODEL DZNR D(BV=10 TBV1=0.75m IS=1E-12 KF=0 RS=0 XTI=0)
.ENDS CUSTOMBLOCK
*
***
*
****** Pinout: OUTA, OUTB, V-, +INB/V+, -INB, -INA, +INA/V+
